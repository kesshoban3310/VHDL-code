Library ieee;
Use ieee.std_logic_1164.all;
ENTITY hex IS
	port(z,y,x,w,z1,y1,x1,w1 : IN STD_LOGIC;
			a,b,c,d,e,f,g,a1,b1,c1,d1,e1,f1,g1      : OUT STD_LOGIC);
end hex;
 
ARCHITECTURE  func OF hex IS 
BEGIN
    a<= (not w and not x and not y and z) or (w and not x and y and z) or (x and not y and not z) or (w and x and not y);
    b<= (w and x and not y and not z) or (not w and x and not y and z) or (w and y and z) or (w and x and y) or (x and y and not z);
    c<= (not w and not x and y and not z) or (w and x and not z) or (w and x and y);
    d<= (not x and not y and z) or (not w and x and not y and not z) or (x and y and z) or (w and not x and y and not z);
    e<= (not w and z) or (not w and x and not y) or (not x and not y and z);
    f<= (not w and not x and z) or (not w and not x and y) or (not w and y and z) or (w and x and not y);
    g<= (not w and not x and not y) or (not w and x and y and z);
    a1<= (not w1 and not x1 and not y1 and z1) or (w1 and not x1 and y1 and z1) or (x1 and not y1 and not z1) or (w1 and x1 and not y1);
    b1<= (w1 and x1 and not y1 and not z1) or (not w1 and x1 and not y1 and z1) or (w1 and y1 and z1) or (w1 and x1 and y1) or (x1 and y1 and not z1);
    c1<= (not w1 and not x1 and y1 and not z1) or (w1 and x1 and not z1) or (w1 and x1 and y1);
    d1<= (not x1 and not y1 and z1) or (not w1 and x1 and not y1 and not z1) or (x1 and y1 and z1) or (w1 and not x1 and y1 and not z1);
    e1<= (not w1 and z1) or (not w1 and x1 and not y1) or (not x1 and not y1 and z1);
    f1<= (not w1 and not x1 and z1) or (not w1 and not x1 and y1) or (not w1 and y1 and z1) or (w1 and x1 and not y1);
    g1<= (not w1 and not x1 and not y1) or (not w1 and x1 and y1 and z1);
END func;